library verilog;
use verilog.vl_types.all;
entity lzw_ctrl is
    generic(
        LIDLE           : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        LINIT_CR        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        WT_LZWST        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        WT_DST1         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        RD_2NDCHAR      : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        WT_DST2         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        \GEN_HASH\      : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WT_HASH         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WT_RHASH        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WR_OREG         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RD_OREG         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RD_OREG2        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHK_CNT         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SP_CHR          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FL_OUT          : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LDONE           : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        done_cr         : out    vl_logic;
        lzw_done        : out    vl_logic;
        gen_hash        : out    vl_logic;
        recal_hash      : out    vl_logic;
        addrb_ioram     : out    vl_logic_vector(11 downto 0);
        enb_ioram       : out    vl_logic;
        web_ioram       : out    vl_logic;
        addrb_outram    : out    vl_logic_vector(11 downto 0);
        enb_outram      : out    vl_logic;
        web_outram      : out    vl_logic;
        addrb_cvram     : out    vl_logic_vector(12 downto 0);
        enb_cvram       : out    vl_logic;
        web_cvram       : out    vl_logic;
        wr_cvdataa      : out    vl_logic_vector(12 downto 0);
        ena_cvram       : out    vl_logic;
        wea_cvram       : out    vl_logic;
        wea_acram       : out    vl_logic;
        wea_pcram       : out    vl_logic;
        write_data      : out    vl_logic;
        read_data       : out    vl_logic;
        write_sp        : out    vl_logic;
        shift_char      : out    vl_logic;
        mux_code_val    : out    vl_logic;
        outram_cnt      : out    vl_logic_vector(11 downto 0);
        init_cr         : in     vl_logic;
        init_lzw        : in     vl_logic;
        char_cnt        : in     vl_logic_vector(11 downto 0);
        not_in_mem      : in     vl_logic;
        in_code_mem     : in     vl_logic;
        match           : in     vl_logic;
        collis          : in     vl_logic;
        valid_dcnt      : in     vl_logic;
        tc_outreg       : in     vl_logic;
        clk             : in     vl_logic;
        rst_n           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LIDLE : constant is 1;
    attribute mti_svvh_generic_type of LINIT_CR : constant is 1;
    attribute mti_svvh_generic_type of WT_LZWST : constant is 1;
    attribute mti_svvh_generic_type of WT_DST1 : constant is 1;
    attribute mti_svvh_generic_type of RD_2NDCHAR : constant is 1;
    attribute mti_svvh_generic_type of WT_DST2 : constant is 1;
    attribute mti_svvh_generic_type of \GEN_HASH\ : constant is 1;
    attribute mti_svvh_generic_type of WT_HASH : constant is 1;
    attribute mti_svvh_generic_type of WT_RHASH : constant is 1;
    attribute mti_svvh_generic_type of WR_OREG : constant is 1;
    attribute mti_svvh_generic_type of RD_OREG : constant is 1;
    attribute mti_svvh_generic_type of RD_OREG2 : constant is 1;
    attribute mti_svvh_generic_type of CHK_CNT : constant is 1;
    attribute mti_svvh_generic_type of SP_CHR : constant is 1;
    attribute mti_svvh_generic_type of FL_OUT : constant is 1;
    attribute mti_svvh_generic_type of LDONE : constant is 1;
end lzw_ctrl;
