library verilog;
use verilog.vl_types.all;
entity test is
end test;
